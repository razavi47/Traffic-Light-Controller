module Seg7dec(x,y); // this module was taken from our Lab 2 submission that we worked on earlier in the semester
	input [3:0] x;
	output [6:0] y;

	assign y[6] = ~x[3]&((~x[2]&~x[1])|(x[2]&x[1]&x[0])) | (x[3]&x[2]&~x[1]&~x[0]);
	assign y[5] = ~x[3]&~x[2]&(x[1] | x[0])|(x[2]&x[0]&(x[3]&~x[1] | ~x[3]&x[1]));
	assign y[4] = ~x[3]&(~x[2]&x[0] | x[2]&~x[1]) | (~x[3]&x[2]&x[1] | x[3]&~x[2]&~x[1])&x[0];
	assign y[3] = (~x[3]&~x[1]&(~x[2]&x[0] | x[2]&~x[0])) | (x[3]&~x[2]&~x[0] | x[2]&x[0])&x[1];
	assign y[2] = ~x[3]&~x[2]&x[1]&~x[0] | x[3]&x[2]&(x[1]|~x[0]);
	assign y[1] = ((~x[3]&x[2]&~x[1] | x[3]&x[1])&x[0]) | ((x[3] | x[1])&(x[2]&~x[0]));
	assign y[0] = (~x[3]&~x[1]&(~x[2]&x[0] | x[2]&~x[0])) | (x[3]&x[0]&(~x[2]&x[1] | x[2]&~x[1]));

endmodule
